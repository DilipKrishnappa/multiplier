package one;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  //`include "design.v"
  //`include "interface.sv"
  `include "transaction.sv"
  `include "sequence.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "scoreboard.sv"
  `include "agent.sv"
  `include "env.sv"
  `include "test.sv"
endpackage
